**********************************************************************
**        Copyright (c) 2014 Carsten Wulff Software, Norway 
** *******************************************************************
** Created       : wulff at 2014-10-2
** Modified      : $Author$ $Date$
** Version       : $Revision$ $HeadURL$
** Description   :  
**********************************************************************


.subckt TGX2_CV A C B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN5 A AVSS AVSS AVSS NCHDL
MN1 B C A AVSS NCHDL
MN2 A C B AVSS NCHDL
MN1b B C A AVSS NCHDL

MP0 AVDD C CN AVSS PCHDL
MP5 A AVDD AVDD AVSS PCHDL
MP1 B CN A AVSS PCHDL
MP2 A CN B AVSS PCHDL
MP1b B CN A AVSS PCHDL

.ends


.SUBCKT PWRSW AVDD_ADC AVDD_CORE AVDD_INT AVSS PWRUP VREF VREF_INT
*.PININFO AVDD_ADC:I AVDD_CORE:I AVSS:I PWRUP:I VREF:I AVDD_INT:O VREF_INT:O

XA1 VREF_INT net011 VREF AVSS  PCHAPL M=31
XB1 AVDD_INT net011 AVDD_ADC AVSS  PCHAPL xoffset=20
XB2 AVDD_INT net011 AVDD_ADC AVSS  PCHAPL  M=30
XC5 VREF_INT AVSS  CAPX20_CV xoffset=20 
XC1 PWRUP net011 AVDD_CORE AVSS  IVX1_CV yoffset=5
XC2 AVSS TAPCELL_CV 
XC2A AVSS TAPCELL_CV 
XC2B AVSS TAPCELL_CV 
XE4 AVDD_INT AVSS  CAPX20_CV 
.ENDS

.SUBCKT MUX8X11 AVDD AVSS D0<11> D0<10> D0<9> D0<8> D0<7> D0<6> 
+ D0<5> D0<4> D0<3> D0<2> D0<1> D0<0> D1<11> D1<10> D1<9> D1<8> D1<7> D1<6> 
+ D1<5> D1<4> D1<3> D1<2> D1<1> D1<0> D2<11> D2<10> D2<9> D2<8> D2<7> D2<6> 
+ D2<5> D2<4> D2<3> D2<2> D2<1> D2<0> D3<11> D3<10> D3<9> D3<8> D3<7> D3<6> 
+ D3<5> D3<4> D3<3> D3<2> D3<1> D3<0> D4<11> D4<10> D4<9> D4<8> D4<7> D4<6> 
+ D4<5> D4<4> D4<3> D4<2> D4<1> D4<0> D5<11> D5<10> D5<9> D5<8> D5<7> D5<6> 
+ D5<5> D5<4> D5<3> D5<2> D5<1> D5<0> D6<11> D6<10> D6<9> D6<8> D6<7> D6<6> 
+ D6<5> D6<4> D6<3> D6<2> D6<1> D6<0> D7<11> D7<10> D7<9> D7<8> D7<7> D7<6> 
+ D7<5> D7<4> D7<3> D7<2> D7<1> D7<0> E S<2> S<1> S<0> Y<11> Y<10> Y<9> Y<8> 
+ Y<7> Y<6> Y<5> Y<4> Y<3> Y<2> Y<1> Y<0>
*.PININFO AVDD:I AVSS:I D0<11>:I D0<10>:I D0<9>:I D0<8>:I D0<7>:I D0<6>:I 
*.PININFO D0<5>:I D0<4>:I D0<3>:I D0<2>:I D0<1>:I D0<0>:I D1<11>:I D1<10>:I 
*.PININFO D1<9>:I D1<8>:I D1<7>:I D1<6>:I D1<5>:I D1<4>:I D1<3>:I D1<2>:I 
*.PININFO D1<1>:I D1<0>:I D2<11>:I D2<10>:I D2<9>:I D2<8>:I D2<7>:I D2<6>:I 
*.PININFO D2<5>:I D2<4>:I D2<3>:I D2<2>:I D2<1>:I D2<0>:I D3<11>:I D3<10>:I 
*.PININFO D3<9>:I D3<8>:I D3<7>:I D3<6>:I D3<5>:I D3<4>:I D3<3>:I D3<2>:I 
*.PININFO D3<1>:I D3<0>:I D4<11>:I D4<10>:I D4<9>:I D4<8>:I D4<7>:I D4<6>:I 
*.PININFO D4<5>:I D4<4>:I D4<3>:I D4<2>:I D4<1>:I D4<0>:I D5<11>:I D5<10>:I 
*.PININFO D5<9>:I D5<8>:I D5<7>:I D5<6>:I D5<5>:I D5<4>:I D5<3>:I D5<2>:I 
*.PININFO D5<1>:I D5<0>:I D6<11>:I D6<10>:I D6<9>:I D6<8>:I D6<7>:I D6<6>:I 
*.PININFO D6<5>:I D6<4>:I D6<3>:I D6<2>:I D6<1>:I D6<0>:I D7<11>:I D7<10>:I 
*.PININFO D7<9>:I D7<8>:I D7<7>:I D7<6>:I D7<5>:I D7<4>:I D7<3>:I D7<2>:I 
*.PININFO D7<1>:I D7<0>:I E:I S<2>:I S<1>:I S<0>:I Y<11>:O Y<10>:O Y<9>:O 
*.PININFO Y<8>:O Y<7>:O Y<6>:O Y<5>:O Y<4>:O Y<3>:O Y<2>:O Y<1>:O Y<0>:O
XA48 D3<11> D3<10> D3<9> D3<8> D3<7> D3<6> D3<5> D3<4> D3<3> D3<2> D3<1> D3<0> 
+ AVDD AVSS T<3> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV 
XB52 D0<11> D0<10> D0<9> D0<8> D0<7> D0<6> D0<5> D0<4> D0<3> D0<2> D0<1> D0<0> 
+ AVDD AVSS T<0> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XC44 D7<11> D7<10> D7<9> D7<8> D7<7> D7<6> D7<5> D7<4> D7<3> D7<2> D7<1> D7<0> 
+ AVDD AVSS T<7> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XD45 D6<11> D6<10> D6<9> D6<8> D6<7> D6<6> D6<5> D6<4> D6<3> D6<2> D6<1> D6<0> 
+ AVDD AVSS T<6> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XE46 D5<11> D5<10> D5<9> D5<8> D5<7> D5<6> D5<5> D5<4> D5<3> D5<2> D5<1> D5<0> 
+ AVDD AVSS T<5> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XF47 D4<11> D4<10> D4<9> D4<8> D4<7> D4<6> D4<5> D4<4> D4<3> D4<2> D4<1> D4<0> 
+ AVDD AVSS T<4> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XG49 D2<11> D2<10> D2<9> D2<8> D2<7> D2<6> D2<5> D2<4> D2<3> D2<2> D2<1> D2<0> 
+ AVDD AVSS T<2> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XH53 D1<11> D1<10> D1<9> D1<8> D1<7> D1<6> D1<5> D1<4> D1<3> D1<2> D1<1> D1<0> 
+ AVDD AVSS T<1> Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> 
+  BUSDRV xoffset=2
XI54 Z<11> Z<10> Z<9> Z<8> Z<7> Z<6> Z<5> Z<4> Z<3> Z<2> Z<1> Z<0> AVDD AVSS E 
+ Y<11> Y<10> Y<9> Y<8> Y<7> Y<6> Y<5> Y<4> Y<3> Y<2> Y<1> Y<0> 
+ DODRV xoffset=6
XJ55  S<2> S<1> S<0> E T<7> T<6> T<5> T<4> T<3> T<2> T<1> T<0> AVDD AVSS 
+ DM3T8X1_CV xoffset=2
.ENDS

.SUBCKT DODRV A<11> A<10> A<9> A<8> A<7> A<6> A<5> A<4> A<3> A<2> 
+ A<1> A<0> AVDD AVSS E Y<11> Y<10> Y<9> Y<8> Y<7> Y<6> Y<5> Y<4> Y<3> Y<2> 
+ Y<1> Y<0>
*.PININFO A<11>:I A<10>:I A<9>:I A<8>:I A<7>:I A<6>:I A<5>:I A<4>:I A<3>:I 
*.PININFO A<2>:I A<1>:I A<0>:I AVDD:I AVSS:I E:I Y<11>:O Y<10>:O Y<9>:O Y<8>:O 
*.PININFO Y<7>:O Y<6>:O Y<5>:O Y<4>:O Y<3>:O Y<2>:O Y<1>:O Y<0>:O

XI5  AVSS  TAPCELL_CV 
XI11 E net17  AVDD AVSS IVX1_CV
XI10<11> A<11>  net17 Y<11> AVDD AVSS NRX1_CV
XI10<10> A<10>  net17 Y<10> AVDD AVSS NRX1_CV
XI10<9> A<9>  net17 Y<9> AVDD AVSS NRX1_CV
XI10<8> A<8>  net17 Y<8> AVDD AVSS NRX1_CV
XI10<7> A<7>  net17 Y<7> AVDD AVSS NRX1_CV
XI10<6> A<6>  net17 Y<6> AVDD AVSS NRX1_CV
XI10<5> A<5>  net17 Y<5> AVDD AVSS NRX1_CV
XI10<4> A<4>  net17 Y<4> AVDD AVSS NRX1_CV
XI10<3> A<3>  net17 Y<3> AVDD AVSS NRX1_CV
XI10<2> A<2>  net17 Y<2> AVDD AVSS NRX1_CV
XI10<1> A<1>  net17 Y<1> AVDD AVSS NRX1_CV
XI10<0> A<0>  net17 Y<0> AVDD AVSS NRX1_CV
.ENDS



.SUBCKT BUSDRV A<11> A<10> A<9> A<8> A<7> A<6> A<5> A<4> A<3> A<2> 
+ A<1> A<0> AVDD AVSS E Y<11> Y<10> Y<9> Y<8> Y<7> Y<6> Y<5> Y<4> Y<3> Y<2> 
+ Y<1> Y<0>
XA2<11> A<11>  E Y<11> AVDD AVSS IVTRICX1_CV
XA2<10> A<10>  E Y<10> AVDD AVSS IVTRICX1_CV
XA2<9> A<9>  E Y<9> AVDD AVSS IVTRICX1_CV
XA2<8> A<8>  E Y<8> AVDD AVSS IVTRICX1_CV
XA2<7> A<7>  E Y<7> AVDD AVSS IVTRICX1_CV
XA2<6> A<6>  E Y<6> AVDD AVSS IVTRICX1_CV
XA2<5> A<5>  E Y<5> AVDD AVSS IVTRICX1_CV
XA2<4> A<4>  E Y<4> AVDD AVSS IVTRICX1_CV
XA2<3> A<3>  E Y<3> AVDD AVSS IVTRICX1_CV
XA2<2> A<2>  E Y<2> AVDD AVSS IVTRICX1_CV
XA2<1> A<1>  E Y<1> AVDD AVSS IVTRICX1_CV
XA2<0> A<0>  E Y<0> AVDD AVSS IVTRICX1_CV
XA4 AVSS TAPCELL_CV
.ENDS



.SUBCKT DI_1V8_ST28N AVDD_1V0 AVDD_1V8 AVSS FROM_PAD_1V8 TO_CORE_1V0
XXC1 FILT_O AVSS  CAPX10_CV angle=180 
XXC2 FROM_PAD_1V8 FILT_O AVSS  RPPO_S0 xoffset=25 yoffset=15

XA5  AVSS  TAPCELL_EV xoffset=20
XA2 FILT_O SCHMITT_O AVDD_1V8 AVSS SCX1_EV

XA5a  AVSS  TAPCELL_EV  yoffset=20
XA3 SCHMITT_O INV_O AVDD_1V0 AVSS  IVX1_EV

XA4 INV_O TO_CORE_1V0 AVDD_1V0 AVSS  IVX8_CV yoffset=15 
XA6  AVSS  TAPCELL_CV 
.ENDS

.SUBCKT SCX1_EV A Y AVDD AVSS
XA2 net10 A AVSS AVSS  NCHDEL 
XA3 sco A net10 AVSS  NCHDEL
XA4a AVDD sco net10 AVSS  NCHDEL
XA4b AVDD sco net10 AVSS  NCHDEL
XA5 Y sco AVSS AVSS  NCHDEL

XB0 net13 A AVDD AVSS  PCHDEL
XB1 sco A net13 AVSS  PCHDEL
XB3a net13 sco AVSS AVSS  PCHDEL
XB3b net13 sco AVSS AVSS  PCHDEL
XB4 Y sco AVDD AVSS  PCHDEL
.ends



.SUBCKT SREGLD8 ARST_N_1V0 AVDD AVSS D<0> PO_1V0<7> PO_1V0<6> 
+ PO_1V0<5> PO_1V0<4> PO_1V0<3> PO_1V0<2> PO_1V0<1> PO_1V0<0> SCK_1V0 SI_1V0 
+ SLOAD_1V0
XI0 AVDD AVSS SCK_1V0 D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> ARST_N_1V0 
+ SI_1V0  SHREG8
XI1  D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> SLOAD_1V0 ARST_N_1V0 PO_1V0<7> 
+ PO_1V0<6> PO_1V0<5> PO_1V0<4> PO_1V0<3> PO_1V0<2> PO_1V0<1> PO_1V0<0> 
+ AVDD AVSS   RGRN8X1_CV
.ENDS


.SUBCKT SHREG8 AVDD AVSS CK D<7> D<6> D<5> D<4> D<3> D<2> D<1> 
+ D<0> RN SI_1V0
XI0 SI_1V0 D<7> D<6> D<5> D<4> D<3> D<2> D<1> CK  RN  D<7> D<6> D<5> D<4> 
+ D<3> D<2> D<1> D<0>  AVDD AVSS  RGRN8X1_CV
.ENDS


.SUBCKT TMX8T1X1_CV A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0>  C<7> C<6> C<5> C<4> C<3> C<2> C<1> C<0> E Y AVDD AVSS

XA12a AVSS TAPCELL_CV
XA12b AVSS TAPCELL_CV
XA12c AVSS TAPCELL_CV
XA12d AVSS TAPCELL_CV
XA12e AVSS TAPCELL_CV
XA20 A<0> C<0> Y_INT AVDD AVSS IVTRICX1_CV
XA12f AVSS TAPCELL_CV
XA12g AVSS TAPCELL_CV
XA12h AVSS TAPCELL_CV
XA21 A<1>  C<1> Y_INT  AVDD AVSS IVTRICX1_CV
XA12i AVSS TAPCELL_CV
XA12j AVSS TAPCELL_CV
XA12k AVSS TAPCELL_CV
XA22 A<2>  C<2> Y_INT  AVDD AVSS IVTRICX1_CV
XA12l AVSS TAPCELL_CV
XA23 A<3>  C<3> Y_INT  AVDD AVSS IVTRICX1_CV

XA12m AVSS TAPCELL_CV
XA12n AVSS TAPCELL_CV
XA10 Y_INT EN Y   AVDD AVSS   NRX1_CV
XA11 E  EN  AVDD AVSS IVX1_CV
XA24 A<4>  C<4> Y_INT  AVDD AVSS IVTRICX1_CV
XA25 A<5>  C<5> Y_INT  AVDD AVSS IVTRICX1_CV
XA12o AVSS TAPCELL_CV
XA12p AVSS TAPCELL_CV
XA12q AVSS TAPCELL_CV
XA12r AVSS TAPCELL_CV
XA12s AVSS TAPCELL_CV
XA12t AVSS TAPCELL_CV
XA12u AVSS TAPCELL_CV
XA12v AVSS TAPCELL_CV

XA26 A<6>  C<6> Y_INT  AVDD AVSS IVTRICX1_CV
XA27 A<7>  C<7> Y_INT AVDD AVSS IVTRICX1_CV
.ENDS

.SUBCKT MUX8T1_CV A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0>  E S<2>  S<1> S<0> Y AVDD AVSS
XB1 A<7> A<6> A<5> A<4> A<3> A<2> A<1> A<0> C<7> C<6> C<5> C<4>  C<3> C<2> C<1> C<0> E Y AVDD AVSS  TMX8T1X1_CV
XA1  S<2> S<1> S<0> E  C<7> C<6> C<5> C<4> C<3> C<2> C<1> C<0>  AVDD AVSS DM3T8X1_CV

.ENDS


************************************************************************
* Library Name: MPW1
* Cell Name:    CKDIV2
* View Name:    schematic
************************************************************************

.SUBCKT CKDIV2 AVDD AVSS CKI CKO CKO50DC RN
XA12v AVSS TAPCELL_CV
XA1 CKI CKIB AVDD AVSS BFX1_CV
XA2 CKIB CKIN AVDD AVSS  IVX1_CV
XA4  QNI CKIN RN CKO50DC QN AVDD AVSS DFRNQNX1_CV
XA3 CKO50DC QNI AVDD AVSS  IVX1_CV
XA5 CKO50DC CKI CKO AVDD AVSS ANX1_CV

.ENDS

.SUBCKT CKDIV256 ARST_N_1V0 AVDD_1V0 AVSS CKO50<7> CKO50<6> 
+ CKO50<5> CKO50<4> CKO50<3> CKO50<2> CKO50<1> CKO50<0> CKO<7> CKO<6> CKO<5> 
+ CKO<4> CKO<3> CKO<2> CKO<1> CKO<0> CK_SQUARE_CV
*.PININFO ARST_N_1V0:I AVDD_1V0:I AVSS:I CK_SQUARE_CV:I CKO50<7>:O CKO50<6>:O 
*.PININFO CKO50<5>:O CKO50<4>:O CKO50<3>:O CKO50<2>:O CKO50<1>:O CKO50<0>:O 
*.PININFO CKO<7>:O CKO<6>:O CKO<5>:O CKO<4>:O CKO<3>:O CKO<2>:O CKO<1>:O 
*.PININFO CKO<0>:O
XA1 AVDD_1V0 AVSS CK_SQUARE_CV CKO<7> CKO50<7> ARST_N_1V0 CKDIV2
XA2 AVDD_1V0 AVSS CKO<7> CKO<6> CKO50<6> ARST_N_1V0  CKDIV2
XB3 AVDD_1V0 AVSS CKO<6> CKO<5> CKO50<5> ARST_N_1V0  CKDIV2
XB4 AVDD_1V0 AVSS CKO<5> CKO<4> CKO50<4> ARST_N_1V0  CKDIV2
XC5 AVDD_1V0 AVSS CKO<4> CKO<3> CKO50<3> ARST_N_1V0  CKDIV2
XC6 AVDD_1V0 AVSS CKO<3> CKO<2> CKO50<2> ARST_N_1V0  CKDIV2
XD7 AVDD_1V0 AVSS CKO<2> CKO<1> CKO50<1> ARST_N_1V0  CKDIV2
XD8 AVDD_1V0 AVSS CKO<1> CKO<0> CKO50<0> ARST_N_1V0  CKDIV2
.ENDS




************************************************************************
* Library Name: MPW1
* Cell Name:    CKGEN
* View Name:    schematic
************************************************************************

.SUBCKT CKGEN ARST_N_1V0 AVDD_1V0 AVSS CK_DIGDIV_1V0<2> 
+ CK_DIGDIV_1V0<1> CK_DIGDIV_1V0<0> CK_DIG_1V0 CK_SAMPLE_1V0 CK_SMPL_1V0<2> 
+ CK_SMPL_1V0<1> CK_SMPL_1V0<0> CK_SQUARE_CV
*.PININFO ARST_N_1V0:I AVDD_1V0:I AVSS:I CK_DIGDIV_1V0<2>:I CK_DIGDIV_1V0<1>:I 
*.PININFO CK_DIGDIV_1V0<0>:I CK_SMPL_1V0<2>:I CK_SMPL_1V0<1>:I 
*.PININFO CK_SMPL_1V0<0>:I CK_SQUARE_CV:I CK_DIG_1V0:O CK_SAMPLE_1V0:O
XI44 net06 AVDD_1V0 AVSS net038 / IVX4_CV
XI46 net011 AVDD_1V0 AVSS net012 / IVX4_CV
XI49 CKO<0> CKO<1> CKO<2> CKO<3> CKO<4> CKO<5> CKO<6> CKO<7> AVDD_1V0 AVSS 
+ net8 CK_SMPL_1V0<2> CK_SMPL_1V0<1> CK_SMPL_1V0<0> net06 / MUX8T1_CV
XI48 CKO50<0> CKO50<1> CKO50<2> CKO50<3> CKO50<4> CKO50<5> CKO50<6> CKO50<7> 
+ AVDD_1V0 AVSS net8 CK_DIGDIV_1V0<2> CK_DIGDIV_1V0<1> CK_DIGDIV_1V0<0> net011 
+ / MUX8T1_CV
XI39 AVDD_1V0 AVSS net8 / TIEH_CV
XI47 net012 AVDD_1V0 AVSS CK_DIG_1V0 / IVX8_CV
XI45 net038 AVDD_1V0 AVSS CK_SAMPLE_1V0 / IVX8_CV
XU1_DIV2<7> AVDD_1V0 AVSS CK_SQUARE_CV CKO<7> CKO50<7> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<6> AVDD_1V0 AVSS CKO<7> CKO<6> CKO50<6> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<5> AVDD_1V0 AVSS CKO<6> CKO<5> CKO50<5> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<4> AVDD_1V0 AVSS CKO<5> CKO<4> CKO50<4> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<3> AVDD_1V0 AVSS CKO<4> CKO<3> CKO50<3> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<2> AVDD_1V0 AVSS CKO<3> CKO<2> CKO50<2> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<1> AVDD_1V0 AVSS CKO<2> CKO<1> CKO50<1> ARST_N_1V0 / 
+ CKDIV2
XU1_DIV2<0> AVDD_1V0 AVSS CKO<1> CKO<0> CKO50<0> ARST_N_1V0 / 
+ CKDIV2
.ENDS

